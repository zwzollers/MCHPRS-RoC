parameter num_outputs = 24;
parameter num_inputs = 16;
parameter num_o_bytes = 8'd3;
parameter num_i_bytes = 8'd3;
parameter input_id_len = 24;
module redstone (tick, inputs, outputs);
        	input tick;
        	input [num_inputs-1:0] inputs;
        	output [num_outputs:0] outputs;

        
    parameter num_outputs = 1, num_inputs = 1;

	wire w107_8_66;
	assign w107_8_66 = inputs[0];
	wire w110_8_66;
	assign w110_8_66 = inputs[1];
	assign outputs[0] = (w108_8_68|w109_8_68);
	wire w114_8_65;
	assign w114_8_65 = inputs[2];
	wire w116_8_127;
	torch #(1'b1) c116_8_127 (.i_clk(tick), .i_in(w118_8_127), .o_out(w116_8_127));
	wire w118_8_127;
	repeater #(1, 1'b0, 0, 0) c118_8_127 (.i_clk(tick), .i_in(w126_8_133), .i_lock(), .o_out(w118_8_127));
	wire w117_8_128;
	torch #(1'b0) c117_8_128 (.i_clk(tick), .i_in(w116_8_127|w117_8_129), .o_out(w117_8_128));
	wire w117_8_129;
	repeater #(1, 1'b0, 0, 0) c117_8_129 (.i_clk(tick), .i_in(w117_8_128), .i_lock(), .o_out(w117_8_129));
	wire w119_8_130;
	torch #(1'b1) c119_8_130 (.i_clk(tick), .i_in(w117_8_128), .o_out(w119_8_130));
	wire w126_8_133;
	repeater #(1, 1'b0, 0, 0) c126_8_133 (.i_clk(tick), .i_in(w126_8_138), .i_lock(), .o_out(w126_8_133));
	wire w117_8_134;
	repeater #(1, 1'b1, 0, 0) c117_8_134 (.i_clk(tick), .i_in(w119_8_130), .i_lock(), .o_out(w117_8_134));
	wire w119_8_135;
	repeater #(1, 1'b1, 1, 0) c119_8_135 (.i_clk(tick), .i_in(w117_8_134), .i_lock(), .o_out(w119_8_135));
	wire w120_8_135;
	repeater #(1, 1'b0, 0, 1) c120_8_135 (.i_clk(tick), .i_in(w121_8_135), .i_lock(w119_8_135), .o_out(w120_8_135));
	wire w121_8_135;
	repeater #(1, 1'b1, 0, 1) c121_8_135 (.i_clk(tick), .i_in(w120_8_135), .i_lock(w119_8_135), .o_out(w121_8_135));
	assign outputs[1] = (w121_8_135);
	wire w126_8_138;
	assign w126_8_138 = inputs[3];
	wire w119_9_133;
	repeater #(1, 1'b0, 0, 0) c119_9_133 (.i_clk(tick), .i_in(w120_8_135), .i_lock(), .o_out(w119_9_133));
	wire w119_10_135;
	repeater #(1, 1'b1, 1, 0) c119_10_135 (.i_clk(tick), .i_in(w117_8_134|w119_9_133), .i_lock(), .o_out(w119_10_135));
	wire w120_10_135;
	repeater #(1, 1'b0, 0, 1) c120_10_135 (.i_clk(tick), .i_in(w121_10_135), .i_lock(w119_10_135), .o_out(w120_10_135));
	wire w121_10_135;
	repeater #(1, 1'b1, 0, 1) c121_10_135 (.i_clk(tick), .i_in(w120_10_135), .i_lock(w122_10_135), .o_out(w121_10_135));
	wire w122_10_135;
	repeater #(1, 1'b1, 1, 0) c122_10_135 (.i_clk(tick), .i_in(w119_9_133|w117_8_134), .i_lock(), .o_out(w122_10_135));
	assign outputs[2] = (w121_10_135);
	wire w119_11_133;
	repeater #(1, 1'b0, 0, 0) c119_11_133 (.i_clk(tick), .i_in(w120_10_135), .i_lock(), .o_out(w119_11_133));
	wire w119_12_135;
	repeater #(1, 1'b1, 1, 0) c119_12_135 (.i_clk(tick), .i_in(w117_8_134|w119_9_133|w119_11_133), .i_lock(), .o_out(w119_12_135));
	wire w120_12_135;
	repeater #(1, 1'b1, 0, 1) c120_12_135 (.i_clk(tick), .i_in(w121_12_135), .i_lock(w119_12_135), .o_out(w120_12_135));
	wire w121_12_135;
	repeater #(1, 1'b0, 0, 1) c121_12_135 (.i_clk(tick), .i_in(w120_12_135), .i_lock(w122_12_135), .o_out(w121_12_135));
	wire w122_12_135;
	repeater #(1, 1'b1, 1, 0) c122_12_135 (.i_clk(tick), .i_in(w119_11_133|w119_9_133|w117_8_134), .i_lock(), .o_out(w122_12_135));
	assign outputs[3] = (w121_12_135);
	wire w119_13_133;
	repeater #(1, 1'b1, 0, 0) c119_13_133 (.i_clk(tick), .i_in(w120_12_135), .i_lock(), .o_out(w119_13_133));
	wire w119_14_135;
	repeater #(1, 1'b1, 1, 0) c119_14_135 (.i_clk(tick), .i_in(w117_8_134|w119_9_133|w119_11_133|w119_13_133), .i_lock(), .o_out(w119_14_135));
	wire w120_14_135;
	repeater #(1, 1'b0, 0, 1) c120_14_135 (.i_clk(tick), .i_in(w121_14_135), .i_lock(w119_14_135), .o_out(w120_14_135));
	wire w121_14_135;
	repeater #(1, 1'b1, 0, 1) c121_14_135 (.i_clk(tick), .i_in(w120_14_135), .i_lock(w122_14_135), .o_out(w121_14_135));
	wire w122_14_135;
	repeater #(1, 1'b1, 1, 0) c122_14_135 (.i_clk(tick), .i_in(w119_13_133|w119_11_133|w119_9_133|w117_8_134), .i_lock(), .o_out(w122_14_135));
	assign outputs[4] = (w121_14_135);
	wire w119_15_133;
	repeater #(1, 1'b0, 0, 0) c119_15_133 (.i_clk(tick), .i_in(w120_14_135), .i_lock(), .o_out(w119_15_133));
	wire w119_16_135;
	repeater #(1, 1'b1, 1, 0) c119_16_135 (.i_clk(tick), .i_in(w117_8_134|w119_9_133|w119_11_133|w119_13_133|w119_15_133), .i_lock(), .o_out(w119_16_135));
	wire w120_16_135;
	repeater #(1, 1'b0, 0, 1) c120_16_135 (.i_clk(tick), .i_in(w121_16_135), .i_lock(w119_16_135), .o_out(w120_16_135));
	wire w121_16_135;
	repeater #(1, 1'b1, 0, 1) c121_16_135 (.i_clk(tick), .i_in(w120_16_135), .i_lock(w122_16_135), .o_out(w121_16_135));
	wire w122_16_135;
	repeater #(1, 1'b1, 1, 0) c122_16_135 (.i_clk(tick), .i_in(w119_15_133|w119_13_133|w119_11_133|w119_9_133|w117_8_134), .i_lock(), .o_out(w122_16_135));
	assign outputs[5] = (w121_16_135);
	wire w119_17_133;
	repeater #(1, 1'b0, 0, 0) c119_17_133 (.i_clk(tick), .i_in(w120_16_135), .i_lock(), .o_out(w119_17_133));
	wire w119_18_135;
	repeater #(1, 1'b1, 1, 0) c119_18_135 (.i_clk(tick), .i_in(w117_8_134|w119_9_133|w119_11_133|w119_13_133|w119_15_133|w119_17_133), .i_lock(), .o_out(w119_18_135));
	wire w120_18_135;
	repeater #(1, 1'b0, 0, 1) c120_18_135 (.i_clk(tick), .i_in(w121_18_135), .i_lock(w119_18_135), .o_out(w120_18_135));
	wire w121_18_135;
	repeater #(1, 1'b1, 0, 1) c121_18_135 (.i_clk(tick), .i_in(w120_18_135), .i_lock(w122_18_135), .o_out(w121_18_135));
	wire w122_18_135;
	repeater #(1, 1'b1, 1, 0) c122_18_135 (.i_clk(tick), .i_in(w119_17_133|w119_15_133|w119_13_133|w119_11_133|w119_9_133|w117_8_134), .i_lock(), .o_out(w122_18_135));
	assign outputs[6] = (w121_18_135);
	wire w119_19_133;
	repeater #(1, 1'b0, 0, 0) c119_19_133 (.i_clk(tick), .i_in(w120_18_135), .i_lock(), .o_out(w119_19_133));
	wire w119_20_135;
	repeater #(1, 1'b1, 1, 0) c119_20_135 (.i_clk(tick), .i_in(w117_8_134|w119_9_133|w119_11_133|w119_13_133|w119_15_133|w119_17_133|w119_19_133), .i_lock(), .o_out(w119_20_135));
	wire w120_20_135;
	repeater #(1, 1'b0, 0, 1) c120_20_135 (.i_clk(tick), .i_in(w121_20_135), .i_lock(w119_20_135), .o_out(w120_20_135));
	wire w121_20_135;
	repeater #(1, 1'b1, 0, 1) c121_20_135 (.i_clk(tick), .i_in(w120_20_135), .i_lock(w122_20_135), .o_out(w121_20_135));
	wire w122_20_135;
	repeater #(1, 1'b1, 1, 0) c122_20_135 (.i_clk(tick), .i_in(w119_19_133|w119_17_133|w119_15_133|w119_13_133|w119_11_133|w119_9_133|w117_8_134), .i_lock(), .o_out(w122_20_135));
	assign outputs[7] = (w121_20_135);
	wire w119_21_133;
	repeater #(1, 1'b0, 0, 0) c119_21_133 (.i_clk(tick), .i_in(w120_20_135), .i_lock(), .o_out(w119_21_133));
	wire w120_22_129;
	torch #(1'b0) c120_22_129 (.i_clk(tick), .i_in(w120_22_132), .o_out(w120_22_129));
	wire w121_22_129;
	repeater #(2, 1'b0, 0, 0) c121_22_129 (.i_clk(tick), .i_in(w120_22_129), .i_lock(), .o_out(w121_22_129));
	wire w121_22_130;
	repeater #(1, 1'b1, 0, 0) c121_22_130 (.i_clk(tick), .i_in(w120_22_132), .i_lock(), .o_out(w121_22_130));
	wire w120_22_132;
	torch #(1'b1) c120_22_132 (.i_clk(tick), .i_in(w120_22_135), .o_out(w120_22_132));
	wire w119_22_135;
	repeater #(1, 1'b1, 1, 0) c119_22_135 (.i_clk(tick), .i_in(w117_8_134|w119_9_133|w119_11_133|w119_13_133|w119_15_133|w119_17_133|w119_19_133|w119_21_133), .i_lock(), .o_out(w119_22_135));
	wire w120_22_135;
	repeater #(1, 1'b0, 0, 1) c120_22_135 (.i_clk(tick), .i_in(w121_22_135), .i_lock(w119_22_135), .o_out(w120_22_135));
	wire w121_22_135;
	repeater #(1, 1'b1, 0, 1) c121_22_135 (.i_clk(tick), .i_in(w120_22_135), .i_lock(w122_22_135), .o_out(w121_22_135));
	wire w122_22_135;
	repeater #(1, 1'b1, 1, 0) c122_22_135 (.i_clk(tick), .i_in(w119_21_133|w119_19_133|w119_17_133|w119_15_133|w119_13_133|w119_11_133|w119_9_133|w117_8_134), .i_lock(), .o_out(w122_22_135));
	assign outputs[8] = (w121_22_135);
	wire w117_24_134;
	repeater #(1, 1'b1, 0, 0) c117_24_134 (.i_clk(tick), .i_in(w121_22_129|w121_22_130), .i_lock(), .o_out(w117_24_134));
	wire w124_24_134;
	repeater #(1, 1'b1, 0, 0) c124_24_134 (.i_clk(tick), .i_in(w121_22_129|w121_22_130), .i_lock(), .o_out(w124_24_134));
	wire w119_24_135;
	repeater #(1, 1'b1, 1, 0) c119_24_135 (.i_clk(tick), .i_in(w117_24_134), .i_lock(), .o_out(w119_24_135));
	wire w120_24_135;
	repeater #(1, 1'b1, 0, 1) c120_24_135 (.i_clk(tick), .i_in(w121_24_135), .i_lock(w119_24_135), .o_out(w120_24_135));
	wire w121_24_135;
	repeater #(1, 1'b0, 0, 1) c121_24_135 (.i_clk(tick), .i_in(w120_24_135), .i_lock(w122_24_135), .o_out(w121_24_135));
	wire w122_24_135;
	repeater #(1, 1'b1, 1, 0) c122_24_135 (.i_clk(tick), .i_in(w124_24_134), .i_lock(), .o_out(w122_24_135));
	assign outputs[9] = (w121_24_135);
	wire w119_25_133;
	repeater #(1, 1'b1, 0, 0) c119_25_133 (.i_clk(tick), .i_in(w120_24_135), .i_lock(), .o_out(w119_25_133));
	wire w119_26_135;
	repeater #(1, 1'b1, 1, 0) c119_26_135 (.i_clk(tick), .i_in(w117_24_134|w119_25_133), .i_lock(), .o_out(w119_26_135));
	wire w120_26_135;
	repeater #(1, 1'b1, 0, 1) c120_26_135 (.i_clk(tick), .i_in(w121_26_135), .i_lock(w119_26_135), .o_out(w120_26_135));
	wire w121_26_135;
	repeater #(1, 1'b0, 0, 1) c121_26_135 (.i_clk(tick), .i_in(w120_26_135), .i_lock(w122_26_135), .o_out(w121_26_135));
	wire w122_26_135;
	repeater #(1, 1'b1, 1, 0) c122_26_135 (.i_clk(tick), .i_in(w119_25_133|w124_24_134), .i_lock(), .o_out(w122_26_135));
	assign outputs[10] = (w121_26_135);
	wire w119_27_133;
	repeater #(1, 1'b1, 0, 0) c119_27_133 (.i_clk(tick), .i_in(w120_26_135), .i_lock(), .o_out(w119_27_133));
	wire w119_28_135;
	repeater #(1, 1'b1, 1, 0) c119_28_135 (.i_clk(tick), .i_in(w117_24_134|w119_25_133|w119_27_133), .i_lock(), .o_out(w119_28_135));
	wire w120_28_135;
	repeater #(1, 1'b1, 0, 1) c120_28_135 (.i_clk(tick), .i_in(w121_28_135), .i_lock(w119_28_135), .o_out(w120_28_135));
	wire w121_28_135;
	repeater #(1, 1'b0, 0, 1) c121_28_135 (.i_clk(tick), .i_in(w120_28_135), .i_lock(w122_28_135), .o_out(w121_28_135));
	wire w122_28_135;
	repeater #(1, 1'b1, 1, 0) c122_28_135 (.i_clk(tick), .i_in(w119_27_133|w119_25_133|w124_24_134), .i_lock(), .o_out(w122_28_135));
	assign outputs[11] = (w121_28_135);
	wire w119_29_133;
	repeater #(1, 1'b1, 0, 0) c119_29_133 (.i_clk(tick), .i_in(w120_28_135), .i_lock(), .o_out(w119_29_133));
	wire w119_30_135;
	repeater #(1, 1'b1, 1, 0) c119_30_135 (.i_clk(tick), .i_in(w117_24_134|w119_25_133|w119_27_133|w119_29_133), .i_lock(), .o_out(w119_30_135));
	wire w120_30_135;
	repeater #(1, 1'b1, 0, 1) c120_30_135 (.i_clk(tick), .i_in(w121_30_135), .i_lock(w119_30_135), .o_out(w120_30_135));
	wire w121_30_135;
	repeater #(1, 1'b0, 0, 1) c121_30_135 (.i_clk(tick), .i_in(w120_30_135), .i_lock(w122_30_135), .o_out(w121_30_135));
	wire w122_30_135;
	repeater #(1, 1'b1, 1, 0) c122_30_135 (.i_clk(tick), .i_in(w119_29_133|w119_27_133|w119_25_133|w124_24_134), .i_lock(), .o_out(w122_30_135));
	assign outputs[12] = (w121_30_135);
	wire w119_31_133;
	repeater #(1, 1'b1, 0, 0) c119_31_133 (.i_clk(tick), .i_in(w120_30_135), .i_lock(), .o_out(w119_31_133));
	wire w119_32_135;
	repeater #(1, 1'b1, 1, 0) c119_32_135 (.i_clk(tick), .i_in(w117_24_134|w119_25_133|w119_27_133|w119_29_133|w119_31_133), .i_lock(), .o_out(w119_32_135));
	wire w120_32_135;
	repeater #(1, 1'b0, 0, 1) c120_32_135 (.i_clk(tick), .i_in(w121_32_135), .i_lock(w119_32_135), .o_out(w120_32_135));
	wire w121_32_135;
	repeater #(1, 1'b1, 0, 1) c121_32_135 (.i_clk(tick), .i_in(w120_32_135), .i_lock(w122_32_135), .o_out(w121_32_135));
	wire w122_32_135;
	repeater #(1, 1'b1, 1, 0) c122_32_135 (.i_clk(tick), .i_in(w119_31_133|w119_29_133|w119_27_133|w119_25_133|w124_24_134), .i_lock(), .o_out(w122_32_135));
	assign outputs[13] = (w121_32_135);
	wire w119_33_133;
	repeater #(1, 1'b0, 0, 0) c119_33_133 (.i_clk(tick), .i_in(w120_32_135), .i_lock(), .o_out(w119_33_133));
	wire w119_34_135;
	repeater #(1, 1'b1, 1, 0) c119_34_135 (.i_clk(tick), .i_in(w117_24_134|w119_25_133|w119_27_133|w119_29_133|w119_31_133|w119_33_133), .i_lock(), .o_out(w119_34_135));
	wire w120_34_135;
	repeater #(1, 1'b1, 0, 1) c120_34_135 (.i_clk(tick), .i_in(w121_34_135), .i_lock(w119_34_135), .o_out(w120_34_135));
	wire w121_34_135;
	repeater #(1, 1'b0, 0, 1) c121_34_135 (.i_clk(tick), .i_in(w120_34_135), .i_lock(w122_34_135), .o_out(w121_34_135));
	wire w122_34_135;
	repeater #(1, 1'b1, 1, 0) c122_34_135 (.i_clk(tick), .i_in(w119_33_133|w119_31_133|w119_29_133|w119_27_133|w119_25_133|w124_24_134), .i_lock(), .o_out(w122_34_135));
	assign outputs[14] = (w121_34_135);
	wire w119_35_133;
	repeater #(1, 1'b1, 0, 0) c119_35_133 (.i_clk(tick), .i_in(w120_34_135), .i_lock(), .o_out(w119_35_133));
	wire w119_36_135;
	repeater #(1, 1'b1, 1, 0) c119_36_135 (.i_clk(tick), .i_in(w117_24_134|w119_25_133|w119_27_133|w119_29_133|w119_31_133|w119_33_133|w119_35_133), .i_lock(), .o_out(w119_36_135));
	wire w120_36_135;
	repeater #(1, 1'b1, 0, 1) c120_36_135 (.i_clk(tick), .i_in(w121_36_135), .i_lock(w119_36_135), .o_out(w120_36_135));
	wire w121_36_135;
	repeater #(1, 1'b0, 0, 1) c121_36_135 (.i_clk(tick), .i_in(w120_36_135), .i_lock(w122_36_135), .o_out(w121_36_135));
	wire w122_36_135;
	repeater #(1, 1'b1, 1, 0) c122_36_135 (.i_clk(tick), .i_in(w119_35_133|w119_33_133|w119_31_133|w119_29_133|w119_27_133|w119_25_133|w124_24_134), .i_lock(), .o_out(w122_36_135));
	assign outputs[15] = (w121_36_135);
	wire w119_37_133;
	repeater #(1, 1'b1, 0, 0) c119_37_133 (.i_clk(tick), .i_in(w120_36_135), .i_lock(), .o_out(w119_37_133));
	wire w120_38_129;
	torch #(1'b0) c120_38_129 (.i_clk(tick), .i_in(w120_38_132), .o_out(w120_38_129));
	wire w121_38_129;
	repeater #(2, 1'b0, 0, 0) c121_38_129 (.i_clk(tick), .i_in(w120_38_129), .i_lock(), .o_out(w121_38_129));
	wire w121_38_130;
	repeater #(1, 1'b1, 0, 0) c121_38_130 (.i_clk(tick), .i_in(w120_38_132), .i_lock(), .o_out(w121_38_130));
	wire w120_38_132;
	torch #(1'b1) c120_38_132 (.i_clk(tick), .i_in(w120_38_135), .o_out(w120_38_132));
	wire w119_38_135;
	repeater #(1, 1'b1, 1, 0) c119_38_135 (.i_clk(tick), .i_in(w117_24_134|w119_25_133|w119_27_133|w119_29_133|w119_31_133|w119_33_133|w119_35_133|w119_37_133), .i_lock(), .o_out(w119_38_135));
	wire w120_38_135;
	repeater #(1, 1'b0, 0, 1) c120_38_135 (.i_clk(tick), .i_in(w121_38_135), .i_lock(w119_38_135), .o_out(w120_38_135));
	wire w121_38_135;
	repeater #(1, 1'b1, 0, 1) c121_38_135 (.i_clk(tick), .i_in(w120_38_135), .i_lock(w122_38_135), .o_out(w121_38_135));
	wire w122_38_135;
	repeater #(1, 1'b1, 1, 0) c122_38_135 (.i_clk(tick), .i_in(w119_37_133|w119_35_133|w119_33_133|w119_31_133|w119_29_133|w119_27_133|w119_25_133|w124_24_134), .i_lock(), .o_out(w122_38_135));
	assign outputs[16] = (w121_38_135);
	wire w117_40_134;
	repeater #(1, 1'b1, 0, 0) c117_40_134 (.i_clk(tick), .i_in(w121_38_129|w121_38_130), .i_lock(), .o_out(w117_40_134));
	wire w124_40_134;
	repeater #(1, 1'b1, 0, 0) c124_40_134 (.i_clk(tick), .i_in(w121_38_129|w121_38_130), .i_lock(), .o_out(w124_40_134));
	wire w119_40_135;
	repeater #(1, 1'b1, 1, 0) c119_40_135 (.i_clk(tick), .i_in(w117_40_134), .i_lock(), .o_out(w119_40_135));
	wire w120_40_135;
	repeater #(1, 1'b0, 0, 1) c120_40_135 (.i_clk(tick), .i_in(w121_40_135), .i_lock(w119_40_135), .o_out(w120_40_135));
	wire w121_40_135;
	repeater #(1, 1'b1, 0, 1) c121_40_135 (.i_clk(tick), .i_in(w120_40_135), .i_lock(w122_40_135), .o_out(w121_40_135));
	wire w122_40_135;
	repeater #(1, 1'b1, 1, 0) c122_40_135 (.i_clk(tick), .i_in(w124_40_134), .i_lock(), .o_out(w122_40_135));
	assign outputs[17] = (w121_40_135);
	wire w119_41_133;
	repeater #(1, 1'b0, 0, 0) c119_41_133 (.i_clk(tick), .i_in(w120_40_135), .i_lock(), .o_out(w119_41_133));
	wire w119_42_135;
	repeater #(1, 1'b1, 1, 0) c119_42_135 (.i_clk(tick), .i_in(w117_40_134|w119_41_133), .i_lock(), .o_out(w119_42_135));
	wire w120_42_135;
	repeater #(1, 1'b1, 0, 1) c120_42_135 (.i_clk(tick), .i_in(w121_42_135), .i_lock(w119_42_135), .o_out(w120_42_135));
	wire w121_42_135;
	repeater #(1, 1'b0, 0, 1) c121_42_135 (.i_clk(tick), .i_in(w120_42_135), .i_lock(w122_42_135), .o_out(w121_42_135));
	wire w122_42_135;
	repeater #(1, 1'b1, 1, 0) c122_42_135 (.i_clk(tick), .i_in(w119_41_133|w124_40_134), .i_lock(), .o_out(w122_42_135));
	assign outputs[18] = (w121_42_135);
	wire w119_43_133;
	repeater #(1, 1'b1, 0, 0) c119_43_133 (.i_clk(tick), .i_in(w120_42_135), .i_lock(), .o_out(w119_43_133));
	wire w119_44_135;
	repeater #(1, 1'b1, 1, 0) c119_44_135 (.i_clk(tick), .i_in(w117_40_134|w119_41_133|w119_43_133), .i_lock(), .o_out(w119_44_135));
	wire w120_44_135;
	repeater #(1, 1'b1, 0, 1) c120_44_135 (.i_clk(tick), .i_in(w121_44_135), .i_lock(w119_44_135), .o_out(w120_44_135));
	wire w121_44_135;
	repeater #(1, 1'b0, 0, 1) c121_44_135 (.i_clk(tick), .i_in(w120_44_135), .i_lock(w122_44_135), .o_out(w121_44_135));
	wire w122_44_135;
	repeater #(1, 1'b1, 1, 0) c122_44_135 (.i_clk(tick), .i_in(w119_43_133|w119_41_133|w124_40_134), .i_lock(), .o_out(w122_44_135));
	assign outputs[19] = (w121_44_135);
	wire w119_45_133;
	repeater #(1, 1'b1, 0, 0) c119_45_133 (.i_clk(tick), .i_in(w120_44_135), .i_lock(), .o_out(w119_45_133));
	wire w119_46_135;
	repeater #(1, 1'b1, 1, 0) c119_46_135 (.i_clk(tick), .i_in(w117_40_134|w119_41_133|w119_43_133|w119_45_133), .i_lock(), .o_out(w119_46_135));
	wire w120_46_135;
	repeater #(1, 1'b0, 0, 1) c120_46_135 (.i_clk(tick), .i_in(w121_46_135), .i_lock(w119_46_135), .o_out(w120_46_135));
	wire w121_46_135;
	repeater #(1, 1'b1, 0, 1) c121_46_135 (.i_clk(tick), .i_in(w120_46_135), .i_lock(w122_46_135), .o_out(w121_46_135));
	wire w122_46_135;
	repeater #(1, 1'b1, 1, 0) c122_46_135 (.i_clk(tick), .i_in(w119_45_133|w119_43_133|w119_41_133|w124_40_134), .i_lock(), .o_out(w122_46_135));
	assign outputs[20] = (w121_46_135);
	wire w119_47_133;
	repeater #(1, 1'b0, 0, 0) c119_47_133 (.i_clk(tick), .i_in(w120_46_135), .i_lock(), .o_out(w119_47_133));
	wire w119_48_135;
	repeater #(1, 1'b1, 1, 0) c119_48_135 (.i_clk(tick), .i_in(w117_40_134|w119_41_133|w119_43_133|w119_45_133|w119_47_133), .i_lock(), .o_out(w119_48_135));
	wire w120_48_135;
	repeater #(1, 1'b1, 0, 1) c120_48_135 (.i_clk(tick), .i_in(w121_48_135), .i_lock(w119_48_135), .o_out(w120_48_135));
	wire w121_48_135;
	repeater #(1, 1'b0, 0, 1) c121_48_135 (.i_clk(tick), .i_in(w120_48_135), .i_lock(w122_48_135), .o_out(w121_48_135));
	wire w122_48_135;
	repeater #(1, 1'b1, 1, 0) c122_48_135 (.i_clk(tick), .i_in(w119_47_133|w119_45_133|w119_43_133|w119_41_133|w124_40_134), .i_lock(), .o_out(w122_48_135));
	assign outputs[21] = (w121_48_135);
	wire w119_49_133;
	repeater #(1, 1'b1, 0, 0) c119_49_133 (.i_clk(tick), .i_in(w120_48_135), .i_lock(), .o_out(w119_49_133));
	wire w119_50_135;
	repeater #(1, 1'b1, 1, 0) c119_50_135 (.i_clk(tick), .i_in(w117_40_134|w119_41_133|w119_43_133|w119_45_133|w119_47_133|w119_49_133), .i_lock(), .o_out(w119_50_135));
	wire w120_50_135;
	repeater #(1, 1'b1, 0, 1) c120_50_135 (.i_clk(tick), .i_in(w121_50_135), .i_lock(w119_50_135), .o_out(w120_50_135));
	wire w121_50_135;
	repeater #(1, 1'b0, 0, 1) c121_50_135 (.i_clk(tick), .i_in(w120_50_135), .i_lock(w122_50_135), .o_out(w121_50_135));
	wire w122_50_135;
	repeater #(1, 1'b1, 1, 0) c122_50_135 (.i_clk(tick), .i_in(w119_49_133|w119_47_133|w119_45_133|w119_43_133|w119_41_133|w124_40_134), .i_lock(), .o_out(w122_50_135));
	assign outputs[22] = (w121_50_135);
	wire w119_51_133;
	repeater #(1, 1'b1, 0, 0) c119_51_133 (.i_clk(tick), .i_in(w120_50_135), .i_lock(), .o_out(w119_51_133));
	wire w119_52_135;
	repeater #(1, 1'b1, 1, 0) c119_52_135 (.i_clk(tick), .i_in(w117_40_134|w119_41_133|w119_43_133|w119_45_133|w119_47_133|w119_49_133|w119_51_133), .i_lock(), .o_out(w119_52_135));
	wire w120_52_135;
	repeater #(1, 1'b1, 0, 1) c120_52_135 (.i_clk(tick), .i_in(w121_52_135), .i_lock(w119_52_135), .o_out(w120_52_135));
	wire w121_52_135;
	repeater #(1, 1'b0, 0, 1) c121_52_135 (.i_clk(tick), .i_in(w120_52_135), .i_lock(w122_52_135), .o_out(w121_52_135));
	wire w122_52_135;
	repeater #(1, 1'b1, 1, 0) c122_52_135 (.i_clk(tick), .i_in(w119_51_133|w119_49_133|w119_47_133|w119_45_133|w119_43_133|w119_41_133|w124_40_134), .i_lock(), .o_out(w122_52_135));
	assign outputs[23] = (w121_52_135);
	wire w119_53_133;
	repeater #(1, 1'b1, 0, 0) c119_53_133 (.i_clk(tick), .i_in(w120_52_135), .i_lock(), .o_out(w119_53_133));
	wire w120_54_129;
	torch #(1'b1) c120_54_129 (.i_clk(tick), .i_in(w120_54_132), .o_out(w120_54_129));
	wire w121_54_129;
	repeater #(2, 1'b1, 0, 0) c121_54_129 (.i_clk(tick), .i_in(w120_54_129), .i_lock(), .o_out(w121_54_129));
	wire w121_54_130;
	repeater #(1, 1'b0, 0, 0) c121_54_130 (.i_clk(tick), .i_in(w120_54_132), .i_lock(), .o_out(w121_54_130));
	wire w120_54_132;
	torch #(1'b0) c120_54_132 (.i_clk(tick), .i_in(w120_54_135), .o_out(w120_54_132));
	wire w119_54_135;
	repeater #(1, 1'b1, 1, 0) c119_54_135 (.i_clk(tick), .i_in(w117_40_134|w119_41_133|w119_43_133|w119_45_133|w119_47_133|w119_49_133|w119_51_133|w119_53_133), .i_lock(), .o_out(w119_54_135));
	wire w120_54_135;
	repeater #(1, 1'b1, 0, 1) c120_54_135 (.i_clk(tick), .i_in(w121_54_135), .i_lock(w119_54_135), .o_out(w120_54_135));
	wire w121_54_135;
	repeater #(1, 1'b0, 0, 1) c121_54_135 (.i_clk(tick), .i_in(w120_54_135), .i_lock(w122_54_135), .o_out(w121_54_135));
	wire w122_54_135;
	repeater #(1, 1'b1, 1, 0) c122_54_135 (.i_clk(tick), .i_in(w119_53_133|w119_51_133|w119_49_133|w119_47_133|w119_45_133|w119_43_133|w119_41_133|w124_40_134), .i_lock(), .o_out(w122_54_135));
	assign outputs[24] = (w121_54_135);
	wire w117_56_134;
	repeater #(1, 1'b1, 0, 0) c117_56_134 (.i_clk(tick), .i_in(w121_54_129|w121_54_130), .i_lock(), .o_out(w117_56_134));
	wire w124_56_134;
	repeater #(1, 1'b1, 0, 0) c124_56_134 (.i_clk(tick), .i_in(w121_54_129|w121_54_130), .i_lock(), .o_out(w124_56_134));
	wire w119_56_135;
	repeater #(1, 1'b1, 1, 0) c119_56_135 (.i_clk(tick), .i_in(w117_56_134), .i_lock(), .o_out(w119_56_135));
	wire w120_56_135;
	repeater #(1, 1'b0, 0, 1) c120_56_135 (.i_clk(tick), .i_in(w121_56_135), .i_lock(w119_56_135), .o_out(w120_56_135));
	wire w121_56_135;
	repeater #(1, 1'b1, 0, 1) c121_56_135 (.i_clk(tick), .i_in(w120_56_135), .i_lock(w122_56_135), .o_out(w121_56_135));
	wire w122_56_135;
	repeater #(1, 1'b1, 1, 0) c122_56_135 (.i_clk(tick), .i_in(w124_56_134), .i_lock(), .o_out(w122_56_135));
	assign outputs[25] = (w121_56_135);
	wire w119_57_133;
	repeater #(1, 1'b0, 0, 0) c119_57_133 (.i_clk(tick), .i_in(w120_56_135), .i_lock(), .o_out(w119_57_133));
	wire w119_58_135;
	repeater #(1, 1'b1, 1, 0) c119_58_135 (.i_clk(tick), .i_in(w117_56_134|w119_57_133), .i_lock(), .o_out(w119_58_135));
	wire w120_58_135;
	repeater #(1, 1'b1, 0, 1) c120_58_135 (.i_clk(tick), .i_in(w121_58_135), .i_lock(w119_58_135), .o_out(w120_58_135));
	wire w121_58_135;
	repeater #(1, 1'b0, 0, 1) c121_58_135 (.i_clk(tick), .i_in(w120_58_135), .i_lock(w122_58_135), .o_out(w121_58_135));
	wire w122_58_135;
	repeater #(1, 1'b1, 1, 0) c122_58_135 (.i_clk(tick), .i_in(w119_57_133|w124_56_134), .i_lock(), .o_out(w122_58_135));
	assign outputs[26] = (w121_58_135);
	wire w119_59_133;
	repeater #(1, 1'b1, 0, 0) c119_59_133 (.i_clk(tick), .i_in(w120_58_135), .i_lock(), .o_out(w119_59_133));
	wire w119_60_135;
	repeater #(1, 1'b1, 1, 0) c119_60_135 (.i_clk(tick), .i_in(w117_56_134|w119_57_133|w119_59_133), .i_lock(), .o_out(w119_60_135));
	wire w120_60_135;
	repeater #(1, 1'b1, 0, 1) c120_60_135 (.i_clk(tick), .i_in(w121_60_135), .i_lock(w119_60_135), .o_out(w120_60_135));
	wire w121_60_135;
	repeater #(1, 1'b0, 0, 1) c121_60_135 (.i_clk(tick), .i_in(w120_60_135), .i_lock(w122_60_135), .o_out(w121_60_135));
	wire w122_60_135;
	repeater #(1, 1'b1, 1, 0) c122_60_135 (.i_clk(tick), .i_in(w119_59_133|w119_57_133|w124_56_134), .i_lock(), .o_out(w122_60_135));
	assign outputs[27] = (w121_60_135);
	wire w119_61_133;
	repeater #(1, 1'b1, 0, 0) c119_61_133 (.i_clk(tick), .i_in(w120_60_135), .i_lock(), .o_out(w119_61_133));
	wire w119_62_135;
	repeater #(1, 1'b1, 1, 0) c119_62_135 (.i_clk(tick), .i_in(w117_56_134|w119_57_133|w119_59_133|w119_61_133), .i_lock(), .o_out(w119_62_135));
	wire w120_62_135;
	repeater #(1, 1'b1, 0, 1) c120_62_135 (.i_clk(tick), .i_in(w121_62_135), .i_lock(w119_62_135), .o_out(w120_62_135));
	wire w121_62_135;
	repeater #(1, 1'b0, 0, 1) c121_62_135 (.i_clk(tick), .i_in(w120_62_135), .i_lock(w122_62_135), .o_out(w121_62_135));
	wire w122_62_135;
	repeater #(1, 1'b1, 1, 0) c122_62_135 (.i_clk(tick), .i_in(w119_61_133|w119_59_133|w119_57_133|w124_56_134), .i_lock(), .o_out(w122_62_135));
	assign outputs[28] = (w121_62_135);
	wire w119_63_133;
	repeater #(1, 1'b1, 0, 0) c119_63_133 (.i_clk(tick), .i_in(w120_62_135), .i_lock(), .o_out(w119_63_133));
	wire w119_64_135;
	repeater #(1, 1'b1, 1, 0) c119_64_135 (.i_clk(tick), .i_in(w117_56_134|w119_57_133|w119_59_133|w119_61_133|w119_63_133), .i_lock(), .o_out(w119_64_135));
	wire w120_64_135;
	repeater #(1, 1'b1, 0, 1) c120_64_135 (.i_clk(tick), .i_in(w121_64_135), .i_lock(w119_64_135), .o_out(w120_64_135));
	wire w121_64_135;
	repeater #(1, 1'b0, 0, 1) c121_64_135 (.i_clk(tick), .i_in(w120_64_135), .i_lock(w122_64_135), .o_out(w121_64_135));
	wire w122_64_135;
	repeater #(1, 1'b1, 1, 0) c122_64_135 (.i_clk(tick), .i_in(w119_63_133|w119_61_133|w119_59_133|w119_57_133|w124_56_134), .i_lock(), .o_out(w122_64_135));
	assign outputs[29] = (w121_64_135);
	wire w119_65_133;
	repeater #(1, 1'b1, 0, 0) c119_65_133 (.i_clk(tick), .i_in(w120_64_135), .i_lock(), .o_out(w119_65_133));
	wire w119_66_135;
	repeater #(1, 1'b1, 1, 0) c119_66_135 (.i_clk(tick), .i_in(w117_56_134|w119_57_133|w119_59_133|w119_61_133|w119_63_133|w119_65_133), .i_lock(), .o_out(w119_66_135));
	wire w120_66_135;
	repeater #(1, 1'b1, 0, 1) c120_66_135 (.i_clk(tick), .i_in(w121_66_135), .i_lock(w119_66_135), .o_out(w120_66_135));
	wire w121_66_135;
	repeater #(1, 1'b0, 0, 1) c121_66_135 (.i_clk(tick), .i_in(w120_66_135), .i_lock(w122_66_135), .o_out(w121_66_135));
	wire w122_66_135;
	repeater #(1, 1'b1, 1, 0) c122_66_135 (.i_clk(tick), .i_in(w119_65_133|w119_63_133|w119_61_133|w119_59_133|w119_57_133|w124_56_134), .i_lock(), .o_out(w122_66_135));
	assign outputs[30] = (w121_66_135);
	wire w119_67_133;
	repeater #(1, 1'b1, 0, 0) c119_67_133 (.i_clk(tick), .i_in(w120_66_135), .i_lock(), .o_out(w119_67_133));
	wire w119_68_135;
	repeater #(1, 1'b1, 1, 0) c119_68_135 (.i_clk(tick), .i_in(w117_56_134|w119_57_133|w119_59_133|w119_61_133|w119_63_133|w119_65_133|w119_67_133), .i_lock(), .o_out(w119_68_135));
	wire w120_68_135;
	repeater #(1, 1'b1, 0, 1) c120_68_135 (.i_clk(tick), .i_in(w121_68_135), .i_lock(w119_68_135), .o_out(w120_68_135));
	wire w121_68_135;
	repeater #(1, 1'b0, 0, 1) c121_68_135 (.i_clk(tick), .i_in(w120_68_135), .i_lock(w122_68_135), .o_out(w121_68_135));
	wire w122_68_135;
	repeater #(1, 1'b1, 1, 0) c122_68_135 (.i_clk(tick), .i_in(w119_67_133|w119_65_133|w119_63_133|w119_61_133|w119_59_133|w119_57_133|w124_56_134), .i_lock(), .o_out(w122_68_135));
	assign outputs[31] = (w121_68_135);
	wire w119_69_133;
	repeater #(1, 1'b1, 0, 0) c119_69_133 (.i_clk(tick), .i_in(w120_68_135), .i_lock(), .o_out(w119_69_133));
	wire w119_70_135;
	repeater #(1, 1'b1, 1, 0) c119_70_135 (.i_clk(tick), .i_in(w117_56_134|w119_57_133|w119_59_133|w119_61_133|w119_63_133|w119_65_133|w119_67_133|w119_69_133), .i_lock(), .o_out(w119_70_135));
	wire w120_70_135;
	repeater #(1, 1'b1, 0, 1) c120_70_135 (.i_clk(tick), .i_in(w121_70_135), .i_lock(w119_70_135), .o_out(w120_70_135));
	wire w121_70_135;
	repeater #(1, 1'b0, 0, 1) c121_70_135 (.i_clk(tick), .i_in(w120_70_135), .i_lock(w122_70_135), .o_out(w121_70_135));
	wire w122_70_135;
	repeater #(1, 1'b1, 1, 0) c122_70_135 (.i_clk(tick), .i_in(w119_69_133|w119_67_133|w119_65_133|w119_63_133|w119_61_133|w119_59_133|w119_57_133|w124_56_134), .i_lock(), .o_out(w122_70_135));
	assign outputs[32] = (w121_70_135);
	wire w128_8_153;
	assign w128_8_153 = inputs[4];
	wire w130_8_153;
	assign w130_8_153 = inputs[5];
	wire w138_8_153;
	assign w138_8_153 = inputs[6];
	wire w140_8_153;
	assign w140_8_153 = inputs[7];
	wire w128_8_156;
	repeater #(1, 1'b0, 0, 0) c128_8_156 (.i_clk(tick), .i_in(w130_8_153|w128_8_153), .i_lock(), .o_out(w128_8_156));
	wire w138_8_156;
	torch #(1'b0) c138_8_156 (.i_clk(tick), .i_in(w139_9_155|w138_9_154), .o_out(w138_8_156));
	assign outputs[33] = (w138_8_156|w140_8_156);
	wire w140_8_156;
	torch #(1'b0) c140_8_156 (.i_clk(tick), .i_in(w139_9_155|w140_9_154), .o_out(w140_8_156));
	assign outputs[34] = (w128_8_156);
	assign outputs[35] = (w128_8_153|w130_8_153);
	wire w134_8_158;
	assign w134_8_158 = inputs[8];
	wire w138_9_154;
	torch #(1'b1) c138_9_154 (.i_clk(tick), .i_in(w138_8_153), .o_out(w138_9_154));
	wire w140_9_154;
	torch #(1'b1) c140_9_154 (.i_clk(tick), .i_in(w140_8_153), .o_out(w140_9_154));
	wire w139_9_155;
	torch #(1'b0) c139_9_155 (.i_clk(tick), .i_in(w138_9_154|w140_9_154), .o_out(w139_9_155));
	wire w148_20_94;
	torch #(1'b1) c148_20_94 (.i_clk(tick), .i_in(w161_26_94|w159_26_94|w157_26_94|w155_26_94), .o_out(w148_20_94));
	wire w158_21_83;
	torch #(1'b0) c158_21_83 (.i_clk(tick), .i_in(w151_24_85), .o_out(w158_21_83));
	wire w154_21_85;
	torch #(1'b0) c154_21_85 (.i_clk(tick), .i_in(w151_23_85), .o_out(w154_21_85));
	wire w151_21_86;
	torch #(1'b1) c151_21_86 (.i_clk(tick), .i_in(w149_23_86), .o_out(w151_21_86));
	wire w154_21_87;
	torch #(1'b0) c154_21_87 (.i_clk(tick), .i_in(w151_23_87), .o_out(w154_21_87));
	wire w147_21_93;
	torch #(1'b0) c147_21_93 (.i_clk(tick), .i_in(w149_22_93), .o_out(w147_21_93));
	wire w148_21_93;
	torch #(1'b0) c148_21_93 (.i_clk(tick), .i_in(w148_20_94), .o_out(w148_21_93));
	wire w154_21_95;
	torch #(1'b0) c154_21_95 (.i_clk(tick), .i_in(w155_22_94), .o_out(w154_21_95));
	wire w156_21_95;
	torch #(1'b0) c156_21_95 (.i_clk(tick), .i_in(w157_22_94), .o_out(w156_21_95));
	wire w149_22_93;
	torch #(1'b1) c149_22_93 (.i_clk(tick), .i_in(w148_21_93), .o_out(w149_22_93));
	wire w155_22_94;
	torch #(1'b1) c155_22_94 (.i_clk(tick), .i_in(w156_25_87|w154_25_83|w154_21_85|w154_21_87|w154_25_87), .o_out(w155_22_94));
	wire w157_22_94;
	torch #(1'b1) c157_22_94 (.i_clk(tick), .i_in(w154_21_85|w156_25_85|w156_25_87|w156_25_89), .o_out(w157_22_94));
	wire w159_22_94;
	torch #(1'b1) c159_22_94 (.i_clk(tick), .i_in(w156_25_89|w154_25_87|w154_21_85|w158_21_83), .o_out(w159_22_94));
	wire w149_22_95;
	torch #(1'b0) c149_22_95 (.i_clk(tick), .i_in(w160_21_95|w158_25_95|w156_21_95|w154_21_95|w150_23_96|w149_21_96), .o_out(w149_22_95));
	wire w149_23_85;
	assign w149_23_85 = inputs[9];
	wire w151_23_85;
	torch #(1'b1) c151_23_85 (.i_clk(tick), .i_in(w149_23_85), .o_out(w151_23_85));
	wire w149_23_86;
	assign w149_23_86 = inputs[10];
	wire w149_23_87;
	assign w149_23_87 = inputs[11];
	wire w151_23_87;
	torch #(1'b1) c151_23_87 (.i_clk(tick), .i_in(w149_23_87), .o_out(w151_23_87));
	wire w155_23_93;
	torch #(1'b1) c155_23_93 (.i_clk(tick), .i_in(w156_25_87|w154_25_83|w154_21_85|w154_21_87|w154_25_87), .o_out(w155_23_93));
	wire w157_23_93;
	torch #(1'b1) c157_23_93 (.i_clk(tick), .i_in(w154_21_85|w156_25_85|w156_25_87|w156_25_89), .o_out(w157_23_93));
	wire w159_23_93;
	torch #(1'b1) c159_23_93 (.i_clk(tick), .i_in(w156_25_89|w154_25_87|w154_21_85|w158_21_83), .o_out(w159_23_93));
	wire w147_23_95;
	torch #(1'b0) c147_23_95 (.i_clk(tick), .i_in(w149_23_96|w147_22_96), .o_out(w147_23_95));
	wire w149_24_85;
	assign w149_24_85 = inputs[12];
	wire w151_24_85;
	torch #(1'b1) c151_24_85 (.i_clk(tick), .i_in(w149_24_85), .o_out(w151_24_85));
	wire w149_24_86;
	assign w149_24_86 = inputs[13];
	wire w151_24_86;
	torch #(1'b1) c151_24_86 (.i_clk(tick), .i_in(w149_24_86), .o_out(w151_24_86));
	wire w149_24_87;
	assign w149_24_87 = inputs[14];
	wire w151_24_87;
	torch #(1'b1) c151_24_87 (.i_clk(tick), .i_in(w149_24_87), .o_out(w151_24_87));
	wire w154_25_83;
	torch #(1'b0) c154_25_83 (.i_clk(tick), .i_in(w151_25_85), .o_out(w154_25_83));
	wire w149_25_85;
	assign w149_25_85 = inputs[15];
	wire w151_25_85;
	torch #(1'b1) c151_25_85 (.i_clk(tick), .i_in(w149_25_85), .o_out(w151_25_85));
	wire w156_25_85;
	torch #(1'b0) c156_25_85 (.i_clk(tick), .i_in(w151_25_86), .o_out(w156_25_85));
	wire w149_25_86;
	assign w149_25_86 = inputs[16];
	wire w151_25_86;
	torch #(1'b1) c151_25_86 (.i_clk(tick), .i_in(w149_25_86), .o_out(w151_25_86));
	wire w149_25_87;
	assign w149_25_87 = inputs[17];
	wire w151_25_87;
	torch #(1'b1) c151_25_87 (.i_clk(tick), .i_in(w149_25_87), .o_out(w151_25_87));
	wire w154_25_87;
	torch #(1'b0) c154_25_87 (.i_clk(tick), .i_in(w151_24_86), .o_out(w154_25_87));
	wire w156_25_87;
	torch #(1'b0) c156_25_87 (.i_clk(tick), .i_in(w151_25_87), .o_out(w156_25_87));
	wire w156_25_89;
	torch #(1'b0) c156_25_89 (.i_clk(tick), .i_in(w151_24_87), .o_out(w156_25_89));
	assign outputs[36] = (w149_22_95|w147_23_95);
	wire w158_25_95;
	torch #(1'b1) c158_25_95 (.i_clk(tick), .i_in(w159_26_94), .o_out(w158_25_95));
	wire w155_26_94;
	torch #(1'b0) c155_26_94 (.i_clk(tick), .i_in(w155_23_93), .o_out(w155_26_94));
	wire w157_26_94;
	torch #(1'b0) c157_26_94 (.i_clk(tick), .i_in(w157_23_93), .o_out(w157_26_94));
	wire w159_26_94;
	torch #(1'b0) c159_26_94 (.i_clk(tick), .i_in(w159_23_93), .o_out(w159_26_94));
	wire w147_20_96;
	torch #(1'b0) c147_20_96 (.i_clk(tick), .i_in(w147_21_93|w148_20_94), .o_out(w147_20_96));
	wire w149_21_96;
	torch #(1'b1) c149_21_96 (.i_clk(tick), .i_in(w147_20_96), .o_out(w149_21_96));
	wire w158_21_97;
	torch #(1'b0) c158_21_97 (.i_clk(tick), .i_in(w159_22_94), .o_out(w158_21_97));
	wire w147_22_96;
	torch #(1'b0) c147_22_96 (.i_clk(tick), .i_in(w149_21_96|w149_22_95), .o_out(w147_22_96));
	wire w149_22_97;
	torch #(1'b0) c149_22_97 (.i_clk(tick), .i_in(w160_21_95|w149_21_96|w156_21_95|w158_21_97|w154_25_97|w150_23_98), .o_out(w149_22_97));
	wire w147_22_98;
	torch #(1'b0) c147_22_98 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_97), .o_out(w147_22_98));
	wire w149_22_99;
	torch #(1'b0) c149_22_99 (.i_clk(tick), .i_in(w160_21_95|w154_25_97|w158_21_97|w149_21_96|w156_21_95|w150_23_100), .o_out(w149_22_99));
	wire w147_22_100;
	torch #(1'b0) c147_22_100 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_99), .o_out(w147_22_100));
	wire w149_22_101;
	torch #(1'b0) c149_22_101 (.i_clk(tick), .i_in(w160_21_95|w158_21_97|w149_21_96|w154_21_95|w156_25_101|w150_23_102), .o_out(w149_22_101));
	wire w147_22_102;
	torch #(1'b0) c147_22_102 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_101), .o_out(w147_22_102));
	wire w149_22_103;
	torch #(1'b0) c149_22_103 (.i_clk(tick), .i_in(w160_21_95|w154_25_97|w149_21_96|w158_25_95|w156_21_95|w150_23_104), .o_out(w149_22_103));
	wire w147_22_104;
	torch #(1'b0) c147_22_104 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_103), .o_out(w147_22_104));
	wire w149_22_105;
	torch #(1'b0) c149_22_105 (.i_clk(tick), .i_in(w160_21_95|w156_25_101|w154_25_97|w158_21_97|w149_21_96|w150_23_106), .o_out(w149_22_105));
	wire w147_22_106;
	torch #(1'b0) c147_22_106 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_105), .o_out(w147_22_106));
	wire w149_22_107;
	torch #(1'b0) c149_22_107 (.i_clk(tick), .i_in(w160_21_95|w156_25_101|w158_21_97|w149_21_96|w154_21_95|w150_23_108), .o_out(w149_22_107));
	wire w147_22_108;
	torch #(1'b0) c147_22_108 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_107), .o_out(w147_22_108));
	wire w149_22_109;
	torch #(1'b0) c149_22_109 (.i_clk(tick), .i_in(w160_21_95|w156_25_101|w154_25_97|w158_21_97|w149_21_96), .o_out(w149_22_109));
	wire w147_22_110;
	torch #(1'b0) c147_22_110 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_109), .o_out(w147_22_110));
	wire w149_23_96;
	torch #(1'b1) c149_23_96 (.i_clk(tick), .i_in(w147_23_95|w149_22_95), .o_out(w149_23_96));
	wire w150_23_96;
	torch #(1'b1) c150_23_96 (.i_clk(tick), .i_in(w147_23_97|w149_22_97), .o_out(w150_23_96));
	wire w147_23_97;
	torch #(1'b0) c147_23_97 (.i_clk(tick), .i_in(w149_23_98|w147_22_98), .o_out(w147_23_97));
	wire w149_23_98;
	torch #(1'b1) c149_23_98 (.i_clk(tick), .i_in(w147_23_97|w149_22_97), .o_out(w149_23_98));
	wire w150_23_98;
	torch #(1'b1) c150_23_98 (.i_clk(tick), .i_in(w147_23_99|w149_22_99), .o_out(w150_23_98));
	wire w147_23_99;
	torch #(1'b0) c147_23_99 (.i_clk(tick), .i_in(w149_23_100|w147_22_100), .o_out(w147_23_99));
	wire w149_23_100;
	torch #(1'b1) c149_23_100 (.i_clk(tick), .i_in(w147_23_99|w149_22_99), .o_out(w149_23_100));
	wire w150_23_100;
	torch #(1'b1) c150_23_100 (.i_clk(tick), .i_in(w147_23_101|w149_22_101), .o_out(w150_23_100));
	wire w147_23_101;
	torch #(1'b0) c147_23_101 (.i_clk(tick), .i_in(w149_23_102|w147_22_102), .o_out(w147_23_101));
	wire w149_23_102;
	torch #(1'b1) c149_23_102 (.i_clk(tick), .i_in(w147_23_101|w149_22_101), .o_out(w149_23_102));
	wire w150_23_102;
	torch #(1'b1) c150_23_102 (.i_clk(tick), .i_in(w147_23_103|w149_22_103), .o_out(w150_23_102));
	wire w147_23_103;
	torch #(1'b0) c147_23_103 (.i_clk(tick), .i_in(w149_23_104|w147_22_104), .o_out(w147_23_103));
	wire w149_23_104;
	torch #(1'b1) c149_23_104 (.i_clk(tick), .i_in(w147_23_103|w149_22_103), .o_out(w149_23_104));
	wire w150_23_104;
	torch #(1'b1) c150_23_104 (.i_clk(tick), .i_in(w147_23_105|w149_22_105), .o_out(w150_23_104));
	wire w147_23_105;
	torch #(1'b0) c147_23_105 (.i_clk(tick), .i_in(w149_23_106|w147_22_106), .o_out(w147_23_105));
	wire w149_23_106;
	torch #(1'b1) c149_23_106 (.i_clk(tick), .i_in(w147_23_105|w149_22_105), .o_out(w149_23_106));
	wire w150_23_106;
	torch #(1'b1) c150_23_106 (.i_clk(tick), .i_in(w147_23_107|w149_22_107), .o_out(w150_23_106));
	wire w147_23_107;
	torch #(1'b0) c147_23_107 (.i_clk(tick), .i_in(w149_23_108|w147_22_108), .o_out(w147_23_107));
	wire w149_23_108;
	torch #(1'b1) c149_23_108 (.i_clk(tick), .i_in(w147_23_107|w149_22_107), .o_out(w149_23_108));
	wire w150_23_108;
	torch #(1'b1) c150_23_108 (.i_clk(tick), .i_in(w147_23_109|w149_22_109), .o_out(w150_23_108));
	wire w147_23_109;
	torch #(1'b0) c147_23_109 (.i_clk(tick), .i_in(w149_23_110|w147_22_110), .o_out(w147_23_109));
	wire w149_23_110;
	torch #(1'b1) c149_23_110 (.i_clk(tick), .i_in(w147_23_109|w149_22_109), .o_out(w149_23_110));
	assign outputs[37] = (w149_22_97|w147_23_97);
	wire w154_25_97;
	torch #(1'b1) c154_25_97 (.i_clk(tick), .i_in(w155_26_94), .o_out(w154_25_97));
	assign outputs[38] = (w149_22_99|w147_23_99);
	assign outputs[39] = (w149_22_101|w147_23_101);
	wire w156_25_101;
	torch #(1'b1) c156_25_101 (.i_clk(tick), .i_in(w157_26_94), .o_out(w156_25_101));
	assign outputs[40] = (w149_22_103|w147_23_103);
	assign outputs[41] = (w149_22_105|w147_23_105);
	assign outputs[42] = (w149_22_107|w147_23_107);
	assign outputs[43] = (w149_22_109|w147_23_109);
	wire w160_21_85;
	torch #(1'b0) c160_21_85 (.i_clk(tick), .i_in(w151_21_86), .o_out(w160_21_85));
	wire w160_21_95;
	torch #(1'b0) c160_21_95 (.i_clk(tick), .i_in(w161_22_94), .o_out(w160_21_95));
	wire w161_22_94;
	torch #(1'b1) c161_22_94 (.i_clk(tick), .i_in(w154_21_87|w160_21_85), .o_out(w161_22_94));
	wire w161_23_93;
	torch #(1'b1) c161_23_93 (.i_clk(tick), .i_in(w154_21_87|w160_21_85), .o_out(w161_23_93));
	wire w161_26_94;
	torch #(1'b0) c161_26_94 (.i_clk(tick), .i_in(w161_23_93), .o_out(w161_26_94));
endmodule
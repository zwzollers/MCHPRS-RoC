module redstone (tick, inputs, outputs);
        	input tick;
        	input [num_inputs-1:0] inputs;
        	output [num_outputs:0] outputs;

        
    parameter num_outputs = 1, num_inputs = 1;

	wire w148_20_94;
	torch #(1'b1) c148_20_94 (.i_clk(tick), .i_in(w161_26_94|w159_26_94|w157_26_94|w155_26_94), .o_out(w148_20_94));
	wire w158_21_83;
	torch #(1'b0) c158_21_83 (.i_clk(tick), .i_in(w151_24_85), .o_out(w158_21_83));
	wire w154_21_85;
	torch #(1'b0) c154_21_85 (.i_clk(tick), .i_in(w151_23_85), .o_out(w154_21_85));
	wire w151_21_86;
	torch #(1'b1) c151_21_86 (.i_clk(tick), .i_in(w149_23_86), .o_out(w151_21_86));
	wire w154_21_87;
	torch #(1'b0) c154_21_87 (.i_clk(tick), .i_in(w151_23_87), .o_out(w154_21_87));
	wire w147_21_93;
	torch #(1'b0) c147_21_93 (.i_clk(tick), .i_in(w149_22_93), .o_out(w147_21_93));
	wire w148_21_93;
	torch #(1'b0) c148_21_93 (.i_clk(tick), .i_in(w148_20_94), .o_out(w148_21_93));
	wire w154_21_95;
	torch #(1'b0) c154_21_95 (.i_clk(tick), .i_in(w155_22_94), .o_out(w154_21_95));
	wire w156_21_95;
	torch #(1'b0) c156_21_95 (.i_clk(tick), .i_in(w157_22_94), .o_out(w156_21_95));
	wire w149_22_93;
	torch #(1'b1) c149_22_93 (.i_clk(tick), .i_in(w148_21_93), .o_out(w149_22_93));
	wire w155_22_94;
	torch #(1'b1) c155_22_94 (.i_clk(tick), .i_in(w156_25_87|w154_25_83|w154_21_85|w154_21_87|w154_25_87), .o_out(w155_22_94));
	wire w157_22_94;
	torch #(1'b1) c157_22_94 (.i_clk(tick), .i_in(w154_21_85|w156_25_85|w156_25_87|w156_25_89), .o_out(w157_22_94));
	wire w159_22_94;
	torch #(1'b1) c159_22_94 (.i_clk(tick), .i_in(w156_25_89|w154_25_87|w154_21_85|w158_21_83), .o_out(w159_22_94));
	wire w149_22_95;
	torch #(1'b0) c149_22_95 (.i_clk(tick), .i_in(w160_21_95|w158_25_95|w156_21_95|w154_21_95|w150_23_96|w149_21_96), .o_out(w149_22_95));
	wire w149_23_85;
	assign w149_23_85 = inputs[0];
	wire w151_23_85;
	torch #(1'b1) c151_23_85 (.i_clk(tick), .i_in(w149_23_85), .o_out(w151_23_85));
	wire w149_23_86;
	assign w149_23_86 = inputs[1];
	wire w149_23_87;
	assign w149_23_87 = inputs[2];
	wire w151_23_87;
	torch #(1'b1) c151_23_87 (.i_clk(tick), .i_in(w149_23_87), .o_out(w151_23_87));
	wire w155_23_93;
	torch #(1'b1) c155_23_93 (.i_clk(tick), .i_in(w156_25_87|w154_25_83|w154_21_85|w154_21_87|w154_25_87), .o_out(w155_23_93));
	wire w157_23_93;
	torch #(1'b1) c157_23_93 (.i_clk(tick), .i_in(w154_21_85|w156_25_85|w156_25_87|w156_25_89), .o_out(w157_23_93));
	wire w159_23_93;
	torch #(1'b1) c159_23_93 (.i_clk(tick), .i_in(w156_25_89|w154_25_87|w154_21_85|w158_21_83), .o_out(w159_23_93));
	wire w147_23_95;
	torch #(1'b0) c147_23_95 (.i_clk(tick), .i_in(w149_23_96|w147_22_96), .o_out(w147_23_95));
	wire w149_24_85;
	assign w149_24_85 = inputs[3];
	wire w151_24_85;
	torch #(1'b1) c151_24_85 (.i_clk(tick), .i_in(w149_24_85), .o_out(w151_24_85));
	wire w149_24_86;
	assign w149_24_86 = inputs[4];
	wire w151_24_86;
	torch #(1'b1) c151_24_86 (.i_clk(tick), .i_in(w149_24_86), .o_out(w151_24_86));
	wire w149_24_87;
	assign w149_24_87 = inputs[5];
	wire w151_24_87;
	torch #(1'b1) c151_24_87 (.i_clk(tick), .i_in(w149_24_87), .o_out(w151_24_87));
	wire w154_25_83;
	torch #(1'b0) c154_25_83 (.i_clk(tick), .i_in(w151_25_85), .o_out(w154_25_83));
	wire w149_25_85;
	assign w149_25_85 = inputs[6];
	wire w151_25_85;
	torch #(1'b1) c151_25_85 (.i_clk(tick), .i_in(w149_25_85), .o_out(w151_25_85));
	wire w156_25_85;
	torch #(1'b0) c156_25_85 (.i_clk(tick), .i_in(w151_25_86), .o_out(w156_25_85));
	wire w149_25_86;
	assign w149_25_86 = inputs[7];
	wire w151_25_86;
	torch #(1'b1) c151_25_86 (.i_clk(tick), .i_in(w149_25_86), .o_out(w151_25_86));
	wire w149_25_87;
	assign w149_25_87 = inputs[8];
	wire w151_25_87;
	torch #(1'b1) c151_25_87 (.i_clk(tick), .i_in(w149_25_87), .o_out(w151_25_87));
	wire w154_25_87;
	torch #(1'b0) c154_25_87 (.i_clk(tick), .i_in(w151_24_86), .o_out(w154_25_87));
	wire w156_25_87;
	torch #(1'b0) c156_25_87 (.i_clk(tick), .i_in(w151_25_87), .o_out(w156_25_87));
	wire w156_25_89;
	torch #(1'b0) c156_25_89 (.i_clk(tick), .i_in(w151_24_87), .o_out(w156_25_89));
	wire w147_25_95;
	assign outputs[0] = (w149_22_95|w147_23_95);
	wire w158_25_95;
	torch #(1'b1) c158_25_95 (.i_clk(tick), .i_in(w159_26_94), .o_out(w158_25_95));
	wire w155_26_94;
	torch #(1'b0) c155_26_94 (.i_clk(tick), .i_in(w155_23_93), .o_out(w155_26_94));
	wire w157_26_94;
	torch #(1'b0) c157_26_94 (.i_clk(tick), .i_in(w157_23_93), .o_out(w157_26_94));
	wire w159_26_94;
	torch #(1'b0) c159_26_94 (.i_clk(tick), .i_in(w159_23_93), .o_out(w159_26_94));
	wire w147_20_96;
	torch #(1'b0) c147_20_96 (.i_clk(tick), .i_in(w147_21_93|w148_20_94), .o_out(w147_20_96));
	wire w149_21_96;
	torch #(1'b1) c149_21_96 (.i_clk(tick), .i_in(w147_20_96), .o_out(w149_21_96));
	wire w158_21_97;
	torch #(1'b0) c158_21_97 (.i_clk(tick), .i_in(w159_22_94), .o_out(w158_21_97));
	wire w147_22_96;
	torch #(1'b0) c147_22_96 (.i_clk(tick), .i_in(w149_21_96|w149_22_95), .o_out(w147_22_96));
	wire w149_22_97;
	torch #(1'b0) c149_22_97 (.i_clk(tick), .i_in(w160_21_95|w149_21_96|w156_21_95|w158_21_97|w154_25_97|w150_23_98), .o_out(w149_22_97));
	wire w147_22_98;
	torch #(1'b0) c147_22_98 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_97), .o_out(w147_22_98));
	wire w149_22_99;
	torch #(1'b0) c149_22_99 (.i_clk(tick), .i_in(w160_21_95|w154_25_97|w158_21_97|w149_21_96|w156_21_95|w150_23_100), .o_out(w149_22_99));
	wire w147_22_100;
	torch #(1'b0) c147_22_100 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_99), .o_out(w147_22_100));
	wire w149_22_101;
	torch #(1'b0) c149_22_101 (.i_clk(tick), .i_in(w160_21_95|w158_21_97|w149_21_96|w154_21_95|w156_25_101|w150_23_102), .o_out(w149_22_101));
	wire w147_22_102;
	torch #(1'b0) c147_22_102 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_101), .o_out(w147_22_102));
	wire w149_22_103;
	torch #(1'b0) c149_22_103 (.i_clk(tick), .i_in(w160_21_95|w154_25_97|w149_21_96|w158_25_95|w156_21_95|w150_23_104), .o_out(w149_22_103));
	wire w147_22_104;
	torch #(1'b0) c147_22_104 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_103), .o_out(w147_22_104));
	wire w149_22_105;
	torch #(1'b0) c149_22_105 (.i_clk(tick), .i_in(w160_21_95|w156_25_101|w154_25_97|w158_21_97|w149_21_96|w150_23_106), .o_out(w149_22_105));
	wire w147_22_106;
	torch #(1'b0) c147_22_106 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_105), .o_out(w147_22_106));
	wire w149_22_107;
	torch #(1'b0) c149_22_107 (.i_clk(tick), .i_in(w160_21_95|w156_25_101|w158_21_97|w149_21_96|w154_21_95|w150_23_108), .o_out(w149_22_107));
	wire w147_22_108;
	torch #(1'b0) c147_22_108 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_107), .o_out(w147_22_108));
	wire w149_22_109;
	torch #(1'b0) c149_22_109 (.i_clk(tick), .i_in(w160_21_95|w156_25_101|w154_25_97|w158_21_97|w149_21_96), .o_out(w149_22_109));
	wire w147_22_110;
	torch #(1'b0) c147_22_110 (.i_clk(tick), .i_in(w149_21_96|w149_21_96|w149_22_109), .o_out(w147_22_110));
	wire w149_23_96;
	torch #(1'b1) c149_23_96 (.i_clk(tick), .i_in(w147_23_95|w149_22_95), .o_out(w149_23_96));
	wire w150_23_96;
	torch #(1'b1) c150_23_96 (.i_clk(tick), .i_in(w147_23_97|w149_22_97), .o_out(w150_23_96));
	wire w147_23_97;
	torch #(1'b0) c147_23_97 (.i_clk(tick), .i_in(w149_23_98|w147_22_98), .o_out(w147_23_97));
	wire w149_23_98;
	torch #(1'b1) c149_23_98 (.i_clk(tick), .i_in(w147_23_97|w149_22_97), .o_out(w149_23_98));
	wire w150_23_98;
	torch #(1'b1) c150_23_98 (.i_clk(tick), .i_in(w147_23_99|w149_22_99), .o_out(w150_23_98));
	wire w147_23_99;
	torch #(1'b0) c147_23_99 (.i_clk(tick), .i_in(w149_23_100|w147_22_100), .o_out(w147_23_99));
	wire w149_23_100;
	torch #(1'b1) c149_23_100 (.i_clk(tick), .i_in(w147_23_99|w149_22_99), .o_out(w149_23_100));
	wire w150_23_100;
	torch #(1'b1) c150_23_100 (.i_clk(tick), .i_in(w147_23_101|w149_22_101), .o_out(w150_23_100));
	wire w147_23_101;
	torch #(1'b0) c147_23_101 (.i_clk(tick), .i_in(w149_23_102|w147_22_102), .o_out(w147_23_101));
	wire w149_23_102;
	torch #(1'b1) c149_23_102 (.i_clk(tick), .i_in(w147_23_101|w149_22_101), .o_out(w149_23_102));
	wire w150_23_102;
	torch #(1'b1) c150_23_102 (.i_clk(tick), .i_in(w147_23_103|w149_22_103), .o_out(w150_23_102));
	wire w147_23_103;
	torch #(1'b0) c147_23_103 (.i_clk(tick), .i_in(w149_23_104|w147_22_104), .o_out(w147_23_103));
	wire w149_23_104;
	torch #(1'b1) c149_23_104 (.i_clk(tick), .i_in(w147_23_103|w149_22_103), .o_out(w149_23_104));
	wire w150_23_104;
	torch #(1'b1) c150_23_104 (.i_clk(tick), .i_in(w147_23_105|w149_22_105), .o_out(w150_23_104));
	wire w147_23_105;
	torch #(1'b0) c147_23_105 (.i_clk(tick), .i_in(w149_23_106|w147_22_106), .o_out(w147_23_105));
	wire w149_23_106;
	torch #(1'b1) c149_23_106 (.i_clk(tick), .i_in(w147_23_105|w149_22_105), .o_out(w149_23_106));
	wire w150_23_106;
	torch #(1'b1) c150_23_106 (.i_clk(tick), .i_in(w147_23_107|w149_22_107), .o_out(w150_23_106));
	wire w147_23_107;
	torch #(1'b0) c147_23_107 (.i_clk(tick), .i_in(w149_23_108|w147_22_108), .o_out(w147_23_107));
	wire w149_23_108;
	torch #(1'b1) c149_23_108 (.i_clk(tick), .i_in(w147_23_107|w149_22_107), .o_out(w149_23_108));
	wire w150_23_108;
	torch #(1'b1) c150_23_108 (.i_clk(tick), .i_in(w147_23_109|w149_22_109), .o_out(w150_23_108));
	wire w147_23_109;
	torch #(1'b0) c147_23_109 (.i_clk(tick), .i_in(w149_23_110|w147_22_110), .o_out(w147_23_109));
	wire w149_23_110;
	torch #(1'b1) c149_23_110 (.i_clk(tick), .i_in(w147_23_109|w149_22_109), .o_out(w149_23_110));
	wire w147_25_97;
	assign outputs[1] = (w149_22_97|w147_23_97);
	wire w154_25_97;
	torch #(1'b1) c154_25_97 (.i_clk(tick), .i_in(w155_26_94), .o_out(w154_25_97));
	wire w147_25_99;
	assign outputs[2] = (w149_22_99|w147_23_99);
	wire w147_25_101;
	assign outputs[3] = (w149_22_101|w147_23_101);
	wire w156_25_101;
	torch #(1'b1) c156_25_101 (.i_clk(tick), .i_in(w157_26_94), .o_out(w156_25_101));
	wire w147_25_103;
	assign outputs[4] = (w149_22_103|w147_23_103);
	wire w147_25_105;
	assign outputs[5] = (w149_22_105|w147_23_105);
	wire w147_25_107;
	assign outputs[6] = (w149_22_107|w147_23_107);
	wire w147_25_109;
	assign outputs[7] = (w149_22_109|w147_23_109);
	wire w160_21_85;
	torch #(1'b0) c160_21_85 (.i_clk(tick), .i_in(w151_21_86), .o_out(w160_21_85));
	wire w160_21_95;
	torch #(1'b0) c160_21_95 (.i_clk(tick), .i_in(w161_22_94), .o_out(w160_21_95));
	wire w161_22_94;
	torch #(1'b1) c161_22_94 (.i_clk(tick), .i_in(w154_21_87|w160_21_85), .o_out(w161_22_94));
	wire w161_23_93;
	torch #(1'b1) c161_23_93 (.i_clk(tick), .i_in(w154_21_87|w160_21_85), .o_out(w161_23_93));
	wire w161_26_94;
	torch #(1'b0) c161_26_94 (.i_clk(tick), .i_in(w161_23_93), .o_out(w161_26_94));
endmodule